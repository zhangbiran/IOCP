class A
{
void hello(int data);
void print(int a, int b);
};

//

//

class B
{
void advanceEquip(int index);
void addBlessValue(int index, A value);
};

class C
{
};